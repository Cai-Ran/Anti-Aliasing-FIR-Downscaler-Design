//support max y decimation factor = 5
module mac_y (
    input clk,
    input rst_n,
    input en_load,
    input [7:0] br1P,
    input [7:0] br2P,
    input [7:0] br3P,
    input [7:0] br4P,
    input [7:0] br5P,
    
    input [1:0] h1_1, h1_2, h1_3,
    input [1:0] h2_1, h2_2, h2_3,
    input [1:0] h3_1, h3_2, h3_3,
    input [1:0] h4_1, h4_2, h4_3,
    input [1:0] h5_1, h5_2, h5_3,

    input [2:0] h1_shft_dir,
    input [2:0] h2_shft_dir,
    input [2:0] h3_shft_dir,
    input [2:0] h4_shft_dir,
    input [2:0] h5_shft_dir,

    input [2:0] normalize,
    output reg en_yout,
    output reg [7:0] out_p
);
    
    reg [7:0] p1, p2, p3, p4, p5;

    //demux
    always @(posedge clk, negedge rst_n) begin
        if (!rst_n)
            {p1, p2, p3, p4, p5} <= 40'b0;
        else if (en_load) begin
            p1 <= br1P;
            p2 <= br2P;
            p3 <= br3P;
            p4 <= br4P;
            p5 <= br5P;
        end
    end

    //barrel shifter
    wire [10:0] h1_1_mul, h1_2_mul, h1_3_mul;
    wire [10:0] h2_1_mul, h2_2_mul, h2_3_mul;
    wire [10:0] h3_1_mul, h3_2_mul, h3_3_mul;
    wire [10:0] h4_1_mul, h4_2_mul, h4_3_mul;
    wire [10:0] h5_1_mul, h5_2_mul, h5_3_mul;
    
    wire [12:0] p1_mul, p2_mul, p3_mul, p4_mul, p5_mul;

    assign h1_1_mul = (!h1_shft_dir[0] && h1_1==0) ? 0 : ((h1_shft_dir[0]) ? p1<<h1_1 : p1>>h1_1);
    assign h1_2_mul = (!h1_shft_dir[1] && h1_2==0) ? 0 : ((h1_shft_dir[1]) ? p1<<h1_2 : p1>>h1_2);
    assign h1_3_mul = (!h1_shft_dir[2] && h1_3==0) ? 0 : ((h1_shft_dir[2]) ? p1<<h1_3 : p1>>h1_3);
    assign p1_mul = h1_1_mul + h1_2_mul + h1_3_mul;

    assign h2_1_mul = (!h2_shft_dir[0] && h2_1==0) ? 0 : ((h2_shft_dir[0]) ? p2 << h2_1 : p2 >> h2_1);
    assign h2_2_mul = (!h2_shft_dir[1] && h2_2==0) ? 0 : ((h2_shft_dir[1]) ? p2 << h2_2 : p2 >> h2_2);
    assign h2_3_mul = (!h2_shft_dir[2] && h2_3==0) ? 0 : ((h2_shft_dir[2]) ? p2 << h2_3 : p2 >> h2_3);
    assign p2_mul = h2_1_mul + h2_2_mul + h2_3_mul;

    assign h3_1_mul = (!h3_shft_dir[0] && h3_1==0) ? 0 : ((h3_shft_dir[0]) ? p3 << h3_1 : p3 >> h3_1);
    assign h3_2_mul = (!h3_shft_dir[1] && h3_2==0) ? 0 : ((h3_shft_dir[1]) ? p3 << h3_2 : p3 >> h3_2);
    assign h3_3_mul = (!h3_shft_dir[2] && h3_3==0) ? 0 : ((h3_shft_dir[2]) ? p3 << h3_3 : p3 >> h3_3);
    assign p3_mul = h3_1_mul + h3_2_mul + h3_3_mul;

    assign h4_1_mul = (!h4_shft_dir[0] && h4_1==0) ? 0 : ((h4_shft_dir[0]) ? p4 << h4_1 : p4 >> h4_1);
    assign h4_2_mul = (!h4_shft_dir[1] && h4_2==0) ? 0 : ((h4_shft_dir[1]) ? p4 << h4_2 : p4 >> h4_2);
    assign h4_3_mul = (!h4_shft_dir[2] && h4_3==0) ? 0 : ((h4_shft_dir[2]) ? p4 << h4_3 : p4 >> h4_3);
    assign p4_mul = h4_1_mul + h4_2_mul + h4_3_mul;

    assign h5_1_mul = (!h5_shft_dir[0] && h5_1==0) ? 0 : ((h5_shft_dir[0]) ? p5 << h5_1 : p5 >> h5_1);
    assign h5_2_mul = (!h5_shft_dir[1] && h5_2==0) ? 0 : ((h5_shft_dir[1]) ? p5 << h5_2 : p5 >> h5_2);
    assign h5_3_mul = (!h5_shft_dir[2] && h5_3==0) ? 0 : ((h5_shft_dir[2]) ? p5 << h5_3 : p5 >> h5_3);
    assign p5_mul = h5_1_mul + h5_2_mul + h5_3_mul;

    wire [14:0] acc_sum;
    assign acc_sum = (p1_mul + p2_mul + p3_mul + p4_mul + p5_mul);


    reg tmp_en, en_out;
    always @(posedge clk, negedge rst_n) begin
        if (!rst_n)
            tmp_en <= 0;
        else
            tmp_en <= en_load;
    end

    always @(negedge clk, negedge rst_n) begin
        if (!rst_n) begin
            en_out<= 0;
            en_yout <= 0;
        end
        else begin 
            en_out <= tmp_en;
            en_yout <= en_out;
        end
    end

    always @(posedge clk, negedge rst_n) begin
        if (!rst_n)
            out_p <= 0;
        else if (tmp_en)
            out_p <= (acc_sum>> normalize);
    end

 
endmodule
