//not depends on resolution
`define MAX_X_DECIMATION_FACTOR_LOG2    3       
`define MAX_Y_DECIMATION_FACTOR_LOG2    3       
`define MAX_ROW_LOG2                    11     
`define MAX_COL_LOG2                    10
`define MAX_RES_TARX                    1600
`define X_ROM_LEN                       512
`define Y_ROM_LEN                       512
`define X_ROM_LEN_LOG2                  9       
`define Y_ROM_LEN_LOG2                  9       
`define NUM_RESLUTION_PAIR              64     
`define RESOLUTION_PAIR_LOG2            6
